module cpu (
	input clk,  
	output cpu_write , 
	output cpu_address,
	output cpu_data
);

endmodule 