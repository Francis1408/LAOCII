


module reserve_station();


endmodule